class pkt_proc_with_ext_mem_sequencer extends uvm_sequencer#(pkt_proc_seq_item);
	`uvm_component_utils(pkt_proc_with_ext_mem_sequencer)
	function new(string name="pkt_proc_with_ext_mem_sequencer",uvm_component parent);
		super.new(name,parent);
	endfunction
endclass

